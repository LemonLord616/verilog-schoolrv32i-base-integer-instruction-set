//
//  schoolRISCV - small RISC-V CPU
//
//  Originally based on Sarah L. Harris MIPS CPU
//  & schoolMIPS project.
//
//  Copyright (c) 2017-2020 Stanislav Zhelnio & Aleksandr Romanov.
//
//  Modified in 2024-2025 by Yuri Panchul & Mike Kuskov.
//

`include "sr_cpu.svh"

module sr_cpu
(
    input           clk,            // clock
    input           rst,            // reset

    output  [31:0]  instr_addr,     // instruction memory address
    input   [31:0]  instr_data,     // instruction memory data

    output  [31:0]  data_addr,      // data memory address
    input   [31:0]  data_data,      // data memory data

    output          invalid_instr,

    input   [ 4:0]  debug_reg_addr, // debug access reg address
    output  [31:0]  debug_reg_data  // debug access reg data
);
    // control wires

    wire        aluZero;
    wire        pcSrc;
    wire        regWrite;
    wire        aluSrc;
    wire        wdSrc;
    wire  [3:0] aluControl;

    // instruction decode wires

    wire [ 6:0] cmdOp;
    wire [ 4:0] rd;
    wire [ 2:0] cmdF3;
    wire [ 4:0] rs1;
    wire [ 4:0] rs2;
    wire [ 6:0] cmdF7;
    wire [31:0] immI;
    wire [31:0] immB;
    wire [31:0] immU;

    // program counter

    wire [31:0] pc;
    wire [31:0] pcBranch = pc + immB;
    wire [31:0] pcPlus4  = pc + 32'd4;
    wire [31:0] pcNext   = pcSrc ? pcBranch : pcPlus4;

    register_with_rst pc_r (clk, rst, pcNext, pc);

    // program memory access

    assign instr_addr = pc >> 2;
    wire [31:0] instr = instr_data;

    // instruction decode

    sr_decode id
    (
        .instr      ( instr       ),
        .cmdOp      ( cmdOp       ),
        .rd         ( rd          ),
        .cmdF3      ( cmdF3       ),
        .rs1        ( rs1         ),
        .rs2        ( rs2         ),
        .cmdF7      ( cmdF7       ),
        .immI       ( immI        ),
        .immB       ( immB        ),
        .immU       ( immU        )
    );

    // register file

    wire [31:0] debug_rd;
    wire [31:0] rd1;
    wire [31:0] rd2;
    wire [31:0] wd3;

    sr_register_file rf
    (
        .clk        ( clk            ),
        .a1         ( rs1            ),
        .a2         ( rs2            ),
        .a3         ( rd             ),
        .rd1        ( rd1            ),
        .rd2        ( rd2            ),
        .wd3        ( wd3            ),
        .we3        ( regWrite       ),

        .dbg_addr   ( debug_reg_addr ),
        .dbg_data   ( debug_rd       )
    );

    // alu

    wire [31:0] srcB = aluSrc ? immI : rd2;
    wire [31:0] aluResult;

    sr_alu alu
    (
        .srcA       ( rd1         ),
        .srcB       ( srcB        ),
        .oper       ( aluControl  ),
        .zero       ( aluZero     ),
        .result     ( aluResult   )
    );

    assign wd3 = wdSrc ? immU : aluResult;

    // control

    sr_control sm_control
    (
        .cmdOp         ( cmdOp         ),
        .cmdF3         ( cmdF3         ),
        .cmdF7         ( cmdF7         ),
        .aluZero       ( aluZero       ),
        .pcSrc         ( pcSrc         ),
        .regWrite      ( regWrite      ),
        .aluSrc        ( aluSrc        ),
        .wdSrc         ( wdSrc         ),
        .aluControl    ( aluControl    ),
        .invalid_instr ( invalid_instr )
    );

    // debug register access

    assign debug_reg_data = (debug_reg_addr != '0) ? debug_rd : pc;

endmodule
